import Configuration::*;
import Payloads::*;
import Enumerations::*;

// do branch target parallel here