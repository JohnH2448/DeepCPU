import Configuration::*;
import Payloads::*;
import Enumerations::*;